interface intf(input logic clk);
  logic rst;
  logic [7:0] a,b;
  logic [3:0] sel;
  logic [7:0] result;
endinterface: intf
